// Radix4PLA0.sv
// PLA for 0-th quotient bit selection 

module Radix4PLA0
(
input logic [5 : 0] r6Abs,
input logic [3 : 0] y4,
output logic q0
);

always_comb
begin

case ({r6Abs, y4})
10'b0001010000: q0 = 1'b1;
10'b0001100000: q0 = 1'b1;
10'b0001110000: q0 = 1'b1;
10'b0010000000: q0 = 1'b1;
10'b0010010000: q0 = 1'b1;
10'b0010100000: q0 = 1'b1;
10'b0010110000: q0 = 1'b1;
10'b0011000000: q0 = 1'b1;
10'b0001010001: q0 = 1'b1;
10'b0001100001: q0 = 1'b1;
10'b0001110001: q0 = 1'b1;
10'b0010000001: q0 = 1'b1;
10'b0010010001: q0 = 1'b1;
10'b0010100001: q0 = 1'b1;
10'b0010110001: q0 = 1'b1;
10'b0011000001: q0 = 1'b1;
10'b0011010001: q0 = 1'b1;
10'b0001100010: q0 = 1'b1;
10'b0001110010: q0 = 1'b1;
10'b0010000010: q0 = 1'b1;
10'b0010010010: q0 = 1'b1;
10'b0010100010: q0 = 1'b1;
10'b0010110010: q0 = 1'b1;
10'b0011000010: q0 = 1'b1;
10'b0011010010: q0 = 1'b1;
10'b0011100010: q0 = 1'b1;
10'b0001100011: q0 = 1'b1;
10'b0001110011: q0 = 1'b1;
10'b0010000011: q0 = 1'b1;
10'b0010010011: q0 = 1'b1;
10'b0010100011: q0 = 1'b1;
10'b0010110011: q0 = 1'b1;
10'b0011000011: q0 = 1'b1;
10'b0011010011: q0 = 1'b1;
10'b0011100011: q0 = 1'b1;
10'b0001100100: q0 = 1'b1;
10'b0001110100: q0 = 1'b1;
10'b0010000100: q0 = 1'b1;
10'b0010010100: q0 = 1'b1;
10'b0010100100: q0 = 1'b1;
10'b0010110100: q0 = 1'b1;
10'b0011000100: q0 = 1'b1;
10'b0011010100: q0 = 1'b1;
10'b0011100100: q0 = 1'b1;
10'b0011110100: q0 = 1'b1;
10'b0001100101: q0 = 1'b1;
10'b0001110101: q0 = 1'b1;
10'b0010000101: q0 = 1'b1;
10'b0010010101: q0 = 1'b1;
10'b0010100101: q0 = 1'b1;
10'b0010110101: q0 = 1'b1;
10'b0011000101: q0 = 1'b1;
10'b0011010101: q0 = 1'b1;
10'b0011100101: q0 = 1'b1;
10'b0011110101: q0 = 1'b1;
10'b0100000101: q0 = 1'b1;
10'b0001110110: q0 = 1'b1;
10'b0010000110: q0 = 1'b1;
10'b0010010110: q0 = 1'b1;
10'b0010100110: q0 = 1'b1;
10'b0010110110: q0 = 1'b1;
10'b0011000110: q0 = 1'b1;
10'b0011010110: q0 = 1'b1;
10'b0011100110: q0 = 1'b1;
10'b0011110110: q0 = 1'b1;
10'b0100000110: q0 = 1'b1;
10'b0100010110: q0 = 1'b1;
10'b0001110111: q0 = 1'b1;
10'b0010000111: q0 = 1'b1;
10'b0010010111: q0 = 1'b1;
10'b0010100111: q0 = 1'b1;
10'b0010110111: q0 = 1'b1;
10'b0011000111: q0 = 1'b1;
10'b0011010111: q0 = 1'b1;
10'b0011100111: q0 = 1'b1;
10'b0011110111: q0 = 1'b1;
10'b0100000111: q0 = 1'b1;
10'b0100010111: q0 = 1'b1;
10'b0100100111: q0 = 1'b1;
10'b0001111000: q0 = 1'b1;
10'b0010001000: q0 = 1'b1;
10'b0010011000: q0 = 1'b1;
10'b0010101000: q0 = 1'b1;
10'b0010111000: q0 = 1'b1;
10'b0011001000: q0 = 1'b1;
10'b0011011000: q0 = 1'b1;
10'b0011101000: q0 = 1'b1;
10'b0011111000: q0 = 1'b1;
10'b0100001000: q0 = 1'b1;
10'b0100011000: q0 = 1'b1;
10'b0100101000: q0 = 1'b1;
10'b0100111000: q0 = 1'b1;
10'b0010001001: q0 = 1'b1;
10'b0010011001: q0 = 1'b1;
10'b0010101001: q0 = 1'b1;
10'b0010111001: q0 = 1'b1;
10'b0011001001: q0 = 1'b1;
10'b0011011001: q0 = 1'b1;
10'b0011101001: q0 = 1'b1;
10'b0011111001: q0 = 1'b1;
10'b0100001001: q0 = 1'b1;
10'b0100011001: q0 = 1'b1;
10'b0100101001: q0 = 1'b1;
10'b0100111001: q0 = 1'b1;
10'b0101001001: q0 = 1'b1;
10'b0010001010: q0 = 1'b1;
10'b0010011010: q0 = 1'b1;
10'b0010101010: q0 = 1'b1;
10'b0010111010: q0 = 1'b1;
10'b0011001010: q0 = 1'b1;
10'b0011011010: q0 = 1'b1;
10'b0011101010: q0 = 1'b1;
10'b0011111010: q0 = 1'b1;
10'b0100001010: q0 = 1'b1;
10'b0100011010: q0 = 1'b1;
10'b0100101010: q0 = 1'b1;
10'b0100111010: q0 = 1'b1;
10'b0101001010: q0 = 1'b1;
10'b0010001011: q0 = 1'b1;
10'b0010011011: q0 = 1'b1;
10'b0010101011: q0 = 1'b1;
10'b0010111011: q0 = 1'b1;
10'b0011001011: q0 = 1'b1;
10'b0011011011: q0 = 1'b1;
10'b0011101011: q0 = 1'b1;
10'b0011111011: q0 = 1'b1;
10'b0100001011: q0 = 1'b1;
10'b0100011011: q0 = 1'b1;
10'b0100101011: q0 = 1'b1;
10'b0100111011: q0 = 1'b1;
10'b0101001011: q0 = 1'b1;
10'b0101011011: q0 = 1'b1;
10'b0010011100: q0 = 1'b1;
10'b0010101100: q0 = 1'b1;
10'b0010111100: q0 = 1'b1;
10'b0011001100: q0 = 1'b1;
10'b0011011100: q0 = 1'b1;
10'b0011101100: q0 = 1'b1;
10'b0011111100: q0 = 1'b1;
10'b0100001100: q0 = 1'b1;
10'b0100011100: q0 = 1'b1;
10'b0100101100: q0 = 1'b1;
10'b0100111100: q0 = 1'b1;
10'b0101001100: q0 = 1'b1;
10'b0101011100: q0 = 1'b1;
10'b0101101100: q0 = 1'b1;
10'b0010011101: q0 = 1'b1;
10'b0010101101: q0 = 1'b1;
10'b0010111101: q0 = 1'b1;
10'b0011001101: q0 = 1'b1;
10'b0011011101: q0 = 1'b1;
10'b0011101101: q0 = 1'b1;
10'b0011111101: q0 = 1'b1;
10'b0100001101: q0 = 1'b1;
10'b0100011101: q0 = 1'b1;
10'b0100101101: q0 = 1'b1;
10'b0100111101: q0 = 1'b1;
10'b0101001101: q0 = 1'b1;
10'b0101011101: q0 = 1'b1;
10'b0101101101: q0 = 1'b1;
10'b0101111101: q0 = 1'b1;
10'b0010011110: q0 = 1'b1;
10'b0010101110: q0 = 1'b1;
10'b0010111110: q0 = 1'b1;
10'b0011001110: q0 = 1'b1;
10'b0011011110: q0 = 1'b1;
10'b0011101110: q0 = 1'b1;
10'b0011111110: q0 = 1'b1;
10'b0100001110: q0 = 1'b1;
10'b0100011110: q0 = 1'b1;
10'b0100101110: q0 = 1'b1;
10'b0100111110: q0 = 1'b1;
10'b0101001110: q0 = 1'b1;
10'b0101011110: q0 = 1'b1;
10'b0101101110: q0 = 1'b1;
10'b0101111110: q0 = 1'b1;
10'b0010101111: q0 = 1'b1;
10'b0010111111: q0 = 1'b1;
10'b0011001111: q0 = 1'b1;
10'b0011011111: q0 = 1'b1;
10'b0011101111: q0 = 1'b1;
10'b0011111111: q0 = 1'b1;
10'b0100001111: q0 = 1'b1;
10'b0100011111: q0 = 1'b1;
10'b0100101111: q0 = 1'b1;
10'b0100111111: q0 = 1'b1;
10'b0101001111: q0 = 1'b1;
10'b0101011111: q0 = 1'b1;
10'b0101101111: q0 = 1'b1;
10'b0101111111: q0 = 1'b1;
10'b0110001111: q0 = 1'b1;
default:        q0 = 1'b0;
endcase
end

endmodule